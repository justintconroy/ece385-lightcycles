library ieee;
use ieee.std_logic_1164.ALL;
use ieee.numeric_std.ALL;

--creates an entity HexDriver which process a 4 bit number and
	--convert it to be used by the 7 pins of the 7 segment display.
	--it will be displayed as the Hexadecimal representation of that
	--four bit number.
entity HexDriver is
	port ( In0 : in std_logic_vector(3 downto 0); --4-bit number input
													--to be displayed.

		Out0 : out std_logic_vector(6 downto 0)); --output in the 
													--form of a seven
													--segment display.
end HexDriver;

architecture Behavioral of HexDriver is

begin

--defines what 7 pin output should be based on 4 bit input.
	with In0 select
	Out0 <= "1000000" when "0000",
		"1111001" when "0001",
		"0100100" when "0010",
		"0110000" when "0011",
		"0011001" when "0100",
		"0010010" when "0101",
		"0000010" when "0110",
		"1111000" when "0111",
		"0000000" when "1000",
		"0010000" when "1001",
		"0001000" when "1010",
		"0000011" when "1011",
		"1000110" when "1100",
		"0100001" when "1101",
		"0000110" when "1110",
		"0001110" when "1111",
		"XXXXXXX" when others;

end Behavioral;
